`define MODULE_NAME FP_Mult_Top
`define NO_CE
`define OVERFLOW
`define UNDERFLOW
`define NAN
`define ZERO
